module test();
	
endmodule